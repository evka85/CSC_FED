------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    20:38:00 2016-08-30
-- Module Name:    GEM_TESTS
-- Description:    This module is the entry point for hardware tests e.g. fiber loopback testing with generated data 
------------------------------------------------------------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.csc_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity csc_tests is
    generic(
        g_NUM_GBT_LINKS     : integer;
        g_NUM_OF_OHs        : integer
    );
    port(
        -- reset
        reset_i                     : in  std_logic;
        
        -- TTC
        ttc_clk_i                   : in  t_ttc_clks;        
        ttc_cmds_i                  : in  t_ttc_cmds;
        
        -- Test control
        loopback_gbt_test_en_i      : in std_logic;
        loopback_8b10b_test_en_i    : in std_logic;
        loopback_8b10b_use_trig_i   : in std_logic;
        
        -- 8b10b links
        daq_8b10b_tx_data_arr_o     : out t_gt_8b10b_tx_data_arr(g_NUM_OF_OHs - 1 downto 0);
        daq_8b10b_rx_data_arr_i     : in  t_gt_8b10b_rx_data_arr(g_NUM_OF_OHs - 1 downto 0);
        trig0_8b10b_rx_data_arr_i   : in  t_gt_8b10b_rx_data_arr(g_NUM_OF_OHs - 1 downto 0);
        trig1_8b10b_rx_data_arr_i   : in  t_gt_8b10b_rx_data_arr(g_NUM_OF_OHs - 1 downto 0);
        
        -- GBT links
        gbt_link_ready_i            : in  std_logic_vector(g_NUM_GBT_LINKS - 1 downto 0);
        gbt_tx_data_arr_o           : out t_gbt_frame_array(g_NUM_GBT_LINKS - 1 downto 0);
        gbt_rx_data_arr_i           : in  t_gbt_frame_array(g_NUM_GBT_LINKS - 1 downto 0);
        
        -- IPbus
        ipb_reset_i                 : in  std_logic;
        ipb_clk_i                   : in  std_logic;
        ipb_miso_o                  : out ipb_rbus;
        ipb_mosi_i                  : in  ipb_wbus        
    );
end csc_tests;

architecture Behavioral of csc_tests is

    -- reset
    signal reset_global                     : std_logic;
    signal reset_local                      : std_logic;
    signal reset                            : std_logic;

    -- control
    signal gbt_loop_through_oh              : std_logic;
    
    -- gbt loopback status
    signal gbt_loop_sync_done_arr           : std_logic_vector(g_NUM_GBT_LINKS - 1 downto 0);
    signal gbt_loop_mega_word_cnt_arr       : t_std32_array(g_NUM_GBT_LINKS - 1 downto 0);
    signal gbt_loop_error_cnt_arr           : t_std32_array(g_NUM_GBT_LINKS - 1 downto 0);
    
    -- 8b10b status
    signal all_8b10b_loop_mega_word_cnt_arr : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal daq_8b10b_loop_sync_done_arr     : std_logic_vector(g_NUM_OF_OHs - 1 downto 0);
    signal daq_8b10b_loop_error_cnt_arr     : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal trig0_8b10b_loop_sync_done_arr   : std_logic_vector(g_NUM_OF_OHs - 1 downto 0);
    signal trig0_8b10b_loop_error_cnt_arr   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal trig1_8b10b_loop_sync_done_arr   : std_logic_vector(g_NUM_OF_OHs - 1 downto 0);
    signal trig1_8b10b_loop_error_cnt_arr   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    
    ------ Register signals begin (this section is generated by <csc_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------    

begin

    --== Resets ==--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => ttc_clk_i.clk_40,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    --== GBT loopback test ==--
    
    i_gbt_loopback_tests : for i in 0 to g_NUM_GBT_LINKS - 1 generate
    
        i_gbt_loopback_test_single : entity work.gbt_loopback_test
            port map(
                reset_i          => reset or not loopback_gbt_test_en_i,
                gbt_clk_i        => ttc_clk_i.clk_40,
                gbt_link_ready_i => gbt_link_ready_i(i),
                gbt_tx_data_o    => gbt_tx_data_arr_o(i),
                gbt_rx_data_i    => gbt_rx_data_arr_i(i),
                oh_in_the_loop_i => gbt_loop_through_oh,
                link_sync_done_o => gbt_loop_sync_done_arr(i),
                mega_word_cnt_o  => gbt_loop_mega_word_cnt_arr(i),
                error_cnt_o      => gbt_loop_error_cnt_arr(i)
            );
    
    end generate;

    --== 8b10b loopback test ==--
    
    i_8b10b_loopback_tests : for i in 0 to g_NUM_OF_OHs - 1 generate
    
        i_gbt_loopback_test_single : entity work.gt_8b10b_loopback_test
            port map(
                reset_i                 => reset or not loopback_8b10b_test_en_i,
                link_clk_i              => ttc_clk_i.clk_160,
                daq_tx_data_o           => daq_8b10b_tx_data_arr_o(i),
                daq_rx_data_i           => daq_8b10b_rx_data_arr_i(i),
                trig0_rx_data_i         => trig0_8b10b_rx_data_arr_i(i),
                trig1_rx_data_i         => trig1_8b10b_rx_data_arr_i(i),
                use_trig_links          => loopback_8b10b_use_trig_i,
                mega_word_cnt_o         => all_8b10b_loop_mega_word_cnt_arr(i),
                daq_link_sync_done_o    => daq_8b10b_loop_sync_done_arr(i),
                daq_error_cnt_o         => daq_8b10b_loop_error_cnt_arr(i),
                trig0_link_sync_done_o  => trig0_8b10b_loop_sync_done_arr(i),
                trig0_error_cnt_o       => trig0_8b10b_loop_error_cnt_arr(i),
                trig1_link_sync_done_o  => trig1_8b10b_loop_sync_done_arr(i),
                trig1_error_cnt_o       => trig1_8b10b_loop_error_cnt_arr(i)
            );
    
    end generate;
    
    --===============================================================================================
    -- this section is generated by <csc_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_GEM_TESTS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_GEM_TESTS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_GEM_TESTS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => ttc_clk_i.clk_40,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0000";
    regs_addresses(1)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1000";
    regs_addresses(2)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1010";
    regs_addresses(3)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1011";
    regs_addresses(4)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1012";
    regs_addresses(5)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1020";
    regs_addresses(6)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1021";
    regs_addresses(7)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1022";
    regs_addresses(8)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1030";
    regs_addresses(9)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1031";
    regs_addresses(10)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1032";
    regs_addresses(11)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1040";
    regs_addresses(12)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1041";
    regs_addresses(13)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1042";
    regs_addresses(14)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1050";
    regs_addresses(15)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1051";
    regs_addresses(16)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1052";
    regs_addresses(17)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1060";
    regs_addresses(18)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1061";
    regs_addresses(19)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1062";
    regs_addresses(20)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2010";
    regs_addresses(21)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2011";
    regs_addresses(22)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2012";
    regs_addresses(23)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2013";
    regs_addresses(24)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2014";
    regs_addresses(25)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2020";
    regs_addresses(26)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2021";
    regs_addresses(27)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2022";
    regs_addresses(28)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2023";
    regs_addresses(29)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2024";

    -- Connect read signals
    regs_read_arr(1)(REG_GEM_TESTS_GBT_LOOPBACK_CTRL_LOOP_THROUGH_OH_BIT) <= gbt_loop_through_oh;
    regs_read_arr(2)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(0);
    regs_read_arr(3)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0);
    regs_read_arr(4)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0);
    regs_read_arr(5)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(1);
    regs_read_arr(6)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1);
    regs_read_arr(7)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1);
    regs_read_arr(8)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(2);
    regs_read_arr(9)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2);
    regs_read_arr(10)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2);
    regs_read_arr(11)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(3);
    regs_read_arr(12)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(3);
    regs_read_arr(13)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(3);
    regs_read_arr(14)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(4);
    regs_read_arr(15)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(4);
    regs_read_arr(16)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(4);
    regs_read_arr(17)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(5);
    regs_read_arr(18)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(5);
    regs_read_arr(19)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(5);
    regs_read_arr(20)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(0);
    regs_read_arr(20)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(0);
    regs_read_arr(20)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(0);
    regs_read_arr(21)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(0);
    regs_read_arr(22)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(0);
    regs_read_arr(23)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(0);
    regs_read_arr(24)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(0);
    regs_read_arr(25)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(1);
    regs_read_arr(25)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(1);
    regs_read_arr(25)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(1);
    regs_read_arr(26)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(1);
    regs_read_arr(27)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(1);
    regs_read_arr(28)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(1);
    regs_read_arr(29)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(1);

    -- Connect write signals
    gbt_loop_through_oh <= regs_write_arr(1)(REG_GEM_TESTS_GBT_LOOPBACK_CTRL_LOOP_THROUGH_OH_BIT);

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults
    regs_defaults(1)(REG_GEM_TESTS_GBT_LOOPBACK_CTRL_LOOP_THROUGH_OH_BIT) <= REG_GEM_TESTS_GBT_LOOPBACK_CTRL_LOOP_THROUGH_OH_DEFAULT;

    -- Define writable regs
    regs_writable_arr(1) <= '1';

    --==== Registers end ============================================================================

end Behavioral;
