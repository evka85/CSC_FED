------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    20:38:00 2016-08-30
-- Module Name:    GEM_TESTS
-- Description:    This module is the entry point for hardware tests e.g. fiber loopback testing with generated data 
------------------------------------------------------------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.csc_pkg.all;
use work.ttc_pkg.all;
use work.gth_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity csc_tests is
    port(
        -- reset
        reset_i                     : in  std_logic;
        
        -- TTC
        ttc_clk_i                   : in  t_ttc_clks;        
        ttc_cmds_i                  : in  t_ttc_cmds;
        
        -- GbE link
        gbe_clk_i                   : in  std_logic;
        gbe_tx_data_o               : out t_gt_8b10b_tx_data;
        gbe_test_enable_o           : out std_logic; 
        
        -- IPbus
        ipb_reset_i                 : in  std_logic;
        ipb_clk_i                   : in  std_logic;
        ipb_miso_o                  : out ipb_rbus;
        ipb_mosi_i                  : in  ipb_wbus        
    );
end csc_tests;

architecture Behavioral of csc_tests is

    -- reset
    signal reset_global         : std_logic;
    signal reset_local          : std_logic;
    signal reset                : std_logic;

    -- GbE test
    signal gbe_test_enable      : std_logic;
    signal gbe_user_data        : std_logic_vector(17 downto 0);
    signal gbe_user_data_en     : std_logic;
    signal gbe_send_en          : std_logic;
    
    ------ Register signals begin (this section is generated by <csc_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_TEST_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_TEST_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_TEST_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_TEST_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_TEST_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_TEST_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_TEST_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_TEST_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_TEST_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------    

begin

    --== Resets ==--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => ttc_clk_i.clk_40,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    --== GbE test ==--
    
    gbe_test_enable_o <= gbe_test_enable;
    
    i_gbe_test : entity work.eth_test
        port map(
            reset_i             => reset,
            gbe_clk_i           => gbe_clk_i,
            gbe_tx_data_o       => gbe_tx_data_o,
            user_data_clk_i     => ipb_clk_i,
            user_data_i         => gbe_user_data(15 downto 0),
            user_data_charisk_i => gbe_user_data(17 downto 16),
            user_data_en_i      => gbe_user_data_en,
            send_en_i           => gbe_send_en
        );

    --===============================================================================================
    -- this section is generated by <csc_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_TEST_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_TEST_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_TEST_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => ipb_clk_i,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_TEST_ADDRESS_MSB downto REG_TEST_ADDRESS_LSB) <= x"00";
    regs_addresses(1)(REG_TEST_ADDRESS_MSB downto REG_TEST_ADDRESS_LSB) <= x"10";
    regs_addresses(2)(REG_TEST_ADDRESS_MSB downto REG_TEST_ADDRESS_LSB) <= x"11";
    regs_addresses(3)(REG_TEST_ADDRESS_MSB downto REG_TEST_ADDRESS_LSB) <= x"12";

    -- Connect read signals
    regs_read_arr(1)(REG_TEST_GBE_TEST_ENABLE_BIT) <= gbe_test_enable;

    -- Connect write signals
    gbe_test_enable <= regs_write_arr(1)(REG_TEST_GBE_TEST_ENABLE_BIT);
    gbe_user_data <= regs_write_arr(2)(REG_TEST_GBE_TEST_PUSH_GBE_DATA_MSB downto REG_TEST_GBE_TEST_PUSH_GBE_DATA_LSB);

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);
    gbe_user_data_en <= regs_write_pulse_arr(2);
    gbe_send_en <= regs_write_pulse_arr(3);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults
    regs_defaults(1)(REG_TEST_GBE_TEST_ENABLE_BIT) <= REG_TEST_GBE_TEST_ENABLE_DEFAULT;
    regs_defaults(2)(REG_TEST_GBE_TEST_PUSH_GBE_DATA_MSB downto REG_TEST_GBE_TEST_PUSH_GBE_DATA_LSB) <= REG_TEST_GBE_TEST_PUSH_GBE_DATA_DEFAULT;

    -- Define writable regs
    regs_writable_arr(1) <= '1';
    regs_writable_arr(2) <= '1';

    --==== Registers end ============================================================================

end Behavioral;
