------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    12:22 2016-05-10
-- Module Name:    trigger
-- Description:    This module handles everything related to sbit cluster data (link synchronization, monitoring, local triggering, matching to L1A and reporting data to DAQ)  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.gth_pkg.all;
use work.csc_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity link_monitor is
    generic(
        g_NUM_OF_DMBs : integer
    );
    port(
        -- reset
        reset_i                 : in  std_logic;
        clk_i                   : in  std_logic;

        -- DMB links
        csc_dmb_rx_usrclk_arr_i : in  std_logic_vector(g_NUM_OF_DMBs - 1 downto 0);
        csc_dmb_rx_data_arr_i   : in  t_gt_8b10b_rx_data_arr(g_NUM_OF_DMBs - 1 downto 0);
        csc_dmb_rx_status_arr_i : in  t_gth_rx_status_arr(g_NUM_OF_DMBs - 1 downto 0);

        -- Spy link
        csc_spy_usrclk_i        : in  std_logic;
        csc_spy_rx_data_i       : in  t_gt_8b10b_rx_data;
        csc_spy_rx_status_i     : in  t_gth_rx_status;
        
        -- IPbus
        ipb_reset_i             : in  std_logic;
        ipb_clk_i               : in  std_logic;
        ipb_miso_o              : out ipb_rbus;
        ipb_mosi_i              : in  ipb_wbus
    );
end link_monitor;

architecture link_monitor_arch of link_monitor is
    
    --=== resets ===--
    
    signal reset_global             : std_logic;
    signal reset_local              : std_logic;
    signal reset                    : std_logic;
    
    --=== counters ===--

    signal dmb_mgt_buf_ovf_arr      : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_mgt_buf_unf_arr      : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_not_in_table_arr     : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_disperr_arr          : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_clk_corr_add_arr     : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_clk_corr_drop_arr    : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);

    signal spy_mgt_buf_ovf          : std_logic_vector(15 downto 0);
    signal spy_mgt_buf_unf          : std_logic_vector(15 downto 0);
    signal spy_not_in_table         : std_logic_vector(15 downto 0);
    signal spy_disperr              : std_logic_vector(15 downto 0);
    signal spy_clk_corr_add         : std_logic_vector(15 downto 0);
    signal spy_clk_corr_drop        : std_logic_vector(15 downto 0);

    ------ Register signals begin (this section is generated by <csc_fed_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_LINKS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------
    
begin

    --================================--
    -- Resets  
    --================================--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => clk_i,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    --================================--
    -- DMB link counetrs  
    --================================--
    
    i_dmbs : for i in 0 to g_NUM_OF_DMBs - 1 generate

        -- elastic buffer overflow counter
        i_cnt_dmb_mgt_buf_ovf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => (csc_dmb_rx_status_arr_i(i).rxbufstatus(2)) and (csc_dmb_rx_status_arr_i(i).rxbufstatus(1)) and (not csc_dmb_rx_status_arr_i(i).rxbufstatus(0)), -- 110
                count_o   => dmb_mgt_buf_ovf_arr(i)
            );
    
        -- elastic buffer underflow counter
        i_cnt_dmb_mgt_buf_unf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => (csc_dmb_rx_status_arr_i(i).rxbufstatus(2)) and (not csc_dmb_rx_status_arr_i(i).rxbufstatus(1)) and (csc_dmb_rx_status_arr_i(i).rxbufstatus(0)), -- 101
                count_o   => dmb_mgt_buf_unf_arr(i)
            );
    
        -- clock correction: idle word insertion counter 
        i_cnt_dmb_clk_corr_add : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => csc_dmb_rx_status_arr_i(i).rxclkcorcnt(1) and csc_dmb_rx_status_arr_i(i).rxclkcorcnt(0), -- 11
                count_o   => dmb_clk_corr_add_arr(i)
            );
    
        -- clock correction: idle word drop counter 
        i_cnt_dmb_clk_corr_drop : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => csc_dmb_rx_status_arr_i(i).rxclkcorcnt(1) xor csc_dmb_rx_status_arr_i(i).rxclkcorcnt(0), -- 10 or 01
                count_o   => dmb_clk_corr_drop_arr(i)
            );

        -- not in table error counter
        i_cnt_dmb_not_in_table : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => csc_dmb_rx_data_arr_i(i).rxnotintable(1) or csc_dmb_rx_data_arr_i(i).rxnotintable(0),
                count_o   => dmb_not_in_table_arr(i)
            );

        -- disparity error counter
        i_cnt_dmb_disperr : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => csc_dmb_rx_data_arr_i(i).rxdisperr(1) or csc_dmb_rx_data_arr_i(i).rxdisperr(0),
                count_o   => dmb_disperr_arr(i)
            );
      
    end generate i_dmbs;
    
    --================================--
    -- Spy link counters  
    --================================--

    -- elastic buffer overflow counter
    i_cnt_spy_mgt_buf_ovf : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => (csc_spy_rx_status_i.rxbufstatus(2)) and (csc_spy_rx_status_i.rxbufstatus(1)) and (not csc_spy_rx_status_i.rxbufstatus(0)), -- 110
            count_o   => spy_mgt_buf_ovf
        );

    -- elastic buffer underflow counter
    i_cnt_spy_mgt_buf_unf : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => (csc_spy_rx_status_i.rxbufstatus(2)) and (not csc_spy_rx_status_i.rxbufstatus(1)) and (csc_spy_rx_status_i.rxbufstatus(0)), -- 101
            count_o   => spy_mgt_buf_unf
        );

    -- clock correction: idle word insertion counter 
    i_cnt_spy_clk_corr_add : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => csc_spy_rx_status_i.rxclkcorcnt(1) and csc_spy_rx_status_i.rxclkcorcnt(0), -- 11
            count_o   => spy_clk_corr_add
        );

    -- clock correction: idle word drop counter 
    i_cnt_spy_clk_corr_drop : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => csc_spy_rx_status_i.rxclkcorcnt(1) xor csc_spy_rx_status_i.rxclkcorcnt(0), -- 10 or 01
            count_o   => spy_clk_corr_drop
        );

    -- not in table error counter
    i_cnt_spy_not_in_table : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => csc_spy_rx_data_i.rxnotintable(1) or csc_spy_rx_data_i.rxnotintable(0),
            count_o   => spy_not_in_table
        );

    -- dispersion error counter
    i_cnt_dmb_disperr : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => csc_spy_rx_data_i.rxdisperr(1) or csc_spy_rx_data_i.rxdisperr(0),
            count_o   => spy_disperr
        );
    
    --===============================================================================================
    -- this section is generated by <csc_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_LINKS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_LINKS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_LINKS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clk_i,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"000";
    regs_addresses(1)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"010";
    regs_addresses(2)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"011";
    regs_addresses(3)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"012";
    regs_addresses(4)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"020";
    regs_addresses(5)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"021";
    regs_addresses(6)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"022";
    regs_addresses(7)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"a00";
    regs_addresses(8)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"a01";
    regs_addresses(9)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"a02";

    -- Connect read signals
    regs_read_arr(1)(REG_LINKS_DMB0_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB0_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(0);
    regs_read_arr(1)(REG_LINKS_DMB0_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB0_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(0);
    regs_read_arr(2)(REG_LINKS_DMB0_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB0_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(0);
    regs_read_arr(2)(REG_LINKS_DMB0_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB0_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(0);
    regs_read_arr(3)(REG_LINKS_DMB0_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB0_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(0);
    regs_read_arr(3)(REG_LINKS_DMB0_DISPERR_CNT_MSB downto REG_LINKS_DMB0_DISPERR_CNT_LSB) <= dmb_disperr_arr(0);
    regs_read_arr(4)(REG_LINKS_DMB1_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB1_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(1);
    regs_read_arr(4)(REG_LINKS_DMB1_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB1_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(1);
    regs_read_arr(5)(REG_LINKS_DMB1_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB1_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(1);
    regs_read_arr(5)(REG_LINKS_DMB1_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB1_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(1);
    regs_read_arr(6)(REG_LINKS_DMB1_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB1_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(1);
    regs_read_arr(6)(REG_LINKS_DMB1_DISPERR_CNT_MSB downto REG_LINKS_DMB1_DISPERR_CNT_LSB) <= dmb_disperr_arr(1);
    regs_read_arr(7)(REG_LINKS_SPY_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_SPY_MGT_BUF_OVF_CNT_LSB) <= spy_mgt_buf_ovf;
    regs_read_arr(7)(REG_LINKS_SPY_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_SPY_MGT_BUF_UNF_CNT_LSB) <= spy_mgt_buf_unf;
    regs_read_arr(8)(REG_LINKS_SPY_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_SPY_CLK_CORR_ADD_CNT_LSB) <= spy_clk_corr_add;
    regs_read_arr(8)(REG_LINKS_SPY_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_SPY_CLK_CORR_DROP_CNT_LSB) <= spy_clk_corr_drop;
    regs_read_arr(9)(REG_LINKS_SPY_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_SPY_NOT_IN_TABLE_CNT_LSB) <= spy_not_in_table;
    regs_read_arr(9)(REG_LINKS_SPY_DISPERR_CNT_MSB downto REG_LINKS_SPY_DISPERR_CNT_LSB) <= spy_disperr;

    -- Connect write signals

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults

    -- Define writable regs

    --==== Registers end ============================================================================
    
end link_monitor_arch;

